module AND (
 input A,B,
 output C );

and a1(C,A,B);
endmodule
