module XOR (
 input A,B,
 output Cout);

xor x1(Cout,A,B);

endmodule
