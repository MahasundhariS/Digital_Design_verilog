module NOR (
 input A, B,
 output C);

nor n1(C,A,B);

endmodule
