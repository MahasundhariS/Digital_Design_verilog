module NOT (
 input A,
 output B);

not n1(B,A);

endmodule
