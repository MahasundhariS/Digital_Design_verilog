module NAND (
 input A, B,
 output Cout );
 
nand n1(C,A,B);

endmodule
